hello
std_logic_vector(to_unsigned(127, 8)),
std_logic_vector(to_unsigned(158, 8)),
std_logic_vector(to_unsigned(187, 8)),
std_logic_vector(to_unsigned(212, 8)),
std_logic_vector(to_unsigned(233, 8)),
std_logic_vector(to_unsigned(247, 8)),
std_logic_vector(to_unsigned(253, 8)),
std_logic_vector(to_unsigned(253, 8)),
std_logic_vector(to_unsigned(244, 8)),
std_logic_vector(to_unsigned(229, 8)),
std_logic_vector(to_unsigned(208, 8)),
std_logic_vector(to_unsigned(181, 8)),
std_logic_vector(to_unsigned(152, 8)),
std_logic_vector(to_unsigned(121, 8)),
std_logic_vector(to_unsigned(90, 8)),
std_logic_vector(to_unsigned(62, 8)),
std_logic_vector(to_unsigned(37, 8)),
std_logic_vector(to_unsigned(18, 8)),
std_logic_vector(to_unsigned(5, 8)),
std_logic_vector(to_unsigned(0, 8)),
std_logic_vector(to_unsigned(2, 8)),
std_logic_vector(to_unsigned(12, 8)),
std_logic_vector(to_unsigned(29, 8)),
std_logic_vector(to_unsigned(51, 8)),
std_logic_vector(to_unsigned(78, 8)),
std_logic_vector(to_unsigned(108, 8)),
std_logic_vector(to_unsigned(139, 8)),
std_logic_vector(to_unsigned(170, 8)),
std_logic_vector(to_unsigned(198, 8)),
std_logic_vector(to_unsigned(221, 8)),
std_logic_vector(to_unsigned(239, 8)),
std_logic_vector(to_unsigned(250, 8)),
std_logic_vector(to_unsigned(254, 8)),
std_logic_vector(to_unsigned(250, 8)),
std_logic_vector(to_unsigned(239, 8)),
std_logic_vector(to_unsigned(221, 8)),
std_logic_vector(to_unsigned(198, 8)),
std_logic_vector(to_unsigned(170, 8)),
std_logic_vector(to_unsigned(139, 8)),
std_logic_vector(to_unsigned(108, 8)),
std_logic_vector(to_unsigned(78, 8)),
std_logic_vector(to_unsigned(51, 8)),
std_logic_vector(to_unsigned(29, 8)),
std_logic_vector(to_unsigned(12, 8)),
std_logic_vector(to_unsigned(2, 8)),
std_logic_vector(to_unsigned(0, 8)),
std_logic_vector(to_unsigned(5, 8)),
std_logic_vector(to_unsigned(18, 8)),
std_logic_vector(to_unsigned(37, 8)),
std_logic_vector(to_unsigned(62, 8)),
std_logic_vector(to_unsigned(90, 8)),
std_logic_vector(to_unsigned(121, 8)),
std_logic_vector(to_unsigned(152, 8)),
std_logic_vector(to_unsigned(181, 8)),
std_logic_vector(to_unsigned(208, 8)),
std_logic_vector(to_unsigned(229, 8)),
std_logic_vector(to_unsigned(244, 8)),
std_logic_vector(to_unsigned(253, 8)),
std_logic_vector(to_unsigned(253, 8)),
std_logic_vector(to_unsigned(247, 8)),
std_logic_vector(to_unsigned(233, 8)),
std_logic_vector(to_unsigned(212, 8)),
std_logic_vector(to_unsigned(187, 8)),
std_logic_vector(to_unsigned(158, 8)),
std_logic_vector(to_unsigned(127, 8)),
std_logic_vector(to_unsigned(96, 8)),
std_logic_vector(to_unsigned(67, 8)),
std_logic_vector(to_unsigned(42, 8)),
std_logic_vector(to_unsigned(21, 8)),
std_logic_vector(to_unsigned(7, 8)),
std_logic_vector(to_unsigned(1, 8)),
std_logic_vector(to_unsigned(1, 8)),
std_logic_vector(to_unsigned(10, 8)),
std_logic_vector(to_unsigned(25, 8)),
std_logic_vector(to_unsigned(46, 8)),
std_logic_vector(to_unsigned(73, 8)),
std_logic_vector(to_unsigned(102, 8)),
std_logic_vector(to_unsigned(133, 8)),
std_logic_vector(to_unsigned(164, 8)),
std_logic_vector(to_unsigned(192, 8)),
std_logic_vector(to_unsigned(217, 8)),
std_logic_vector(to_unsigned(236, 8)),
std_logic_vector(to_unsigned(249, 8)),
std_logic_vector(to_unsigned(254, 8)),
std_logic_vector(to_unsigned(252, 8)),
std_logic_vector(to_unsigned(242, 8)),
std_logic_vector(to_unsigned(225, 8)),
std_logic_vector(to_unsigned(203, 8)),
std_logic_vector(to_unsigned(176, 8)),
std_logic_vector(to_unsigned(146, 8)),
std_logic_vector(to_unsigned(115, 8)),
std_logic_vector(to_unsigned(84, 8)),
std_logic_vector(to_unsigned(56, 8)),
std_logic_vector(to_unsigned(33, 8)),
std_logic_vector(to_unsigned(15, 8)),
std_logic_vector(to_unsigned(4, 8)),
std_logic_vector(to_unsigned(0, 8)),
std_logic_vector(to_unsigned(4, 8)),
std_logic_vector(to_unsigned(15, 8)),
std_logic_vector(to_unsigned(33, 8)),
std_logic_vector(to_unsigned(56, 8)),
std_logic_vector(to_unsigned(84, 8)),
std_logic_vector(to_unsigned(115, 8)),
std_logic_vector(to_unsigned(146, 8)),
std_logic_vector(to_unsigned(176, 8)),
std_logic_vector(to_unsigned(203, 8)),
std_logic_vector(to_unsigned(225, 8)),
std_logic_vector(to_unsigned(242, 8)),
std_logic_vector(to_unsigned(252, 8)),
std_logic_vector(to_unsigned(254, 8)),
std_logic_vector(to_unsigned(249, 8)),
std_logic_vector(to_unsigned(236, 8)),
std_logic_vector(to_unsigned(217, 8)),
std_logic_vector(to_unsigned(192, 8)),
std_logic_vector(to_unsigned(164, 8)),
std_logic_vector(to_unsigned(133, 8)),
std_logic_vector(to_unsigned(102, 8)),
std_logic_vector(to_unsigned(73, 8)),
std_logic_vector(to_unsigned(46, 8)),
std_logic_vector(to_unsigned(25, 8)),
std_logic_vector(to_unsigned(10, 8)),
std_logic_vector(to_unsigned(1, 8)),
std_logic_vector(to_unsigned(1, 8)),
std_logic_vector(to_unsigned(7, 8)),
std_logic_vector(to_unsigned(21, 8)),
std_logic_vector(to_unsigned(42, 8)),
std_logic_vector(to_unsigned(67, 8)),
std_logic_vector(to_unsigned(96, 8)),
